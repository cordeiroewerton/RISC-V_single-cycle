module CPU-0.1(); //Definir as entradas

	logic [31:0] w_inst;

endmodule
