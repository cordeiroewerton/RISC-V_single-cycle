module Instr_Mem(input logic[7:0] A, output logic[31:0] RD);
	always_comb begin
		case(A)
			8'h00: RD = 32'b000000000011_00000_000_00001_0010011;
			8'h04: RD = 32'b000000001001_00000_000_00010_0010011;
			8'h08: RD = 32'b0000000_00010_00001_000_00010_0110011;
			8'h0C: RD = 32'b0000000_00010_00001_111_00011_0110011;
			8'h10: RD = 32'b0000000_00010_00001_110_00100_0110011;
			8'h14: RD = 32'b0000000_00100_00011_010_00101_0110011;
			8'h18: RD = 32'b0100000_00101_00100_000_00110_0110011;
			default: RD = 32'b000000_00000_00000_00000_00000_000000;
		endcase
	end
endmodule 
