module Instr_Mem(input logic[7:0] A, output logic[31:0] RD);
	always_comb begin
		case(A)
			8'h00: RD = 32'b00001010101100000000000010010011;
			8'h04: RD = 32'b00000000000100000000010100100011;
			8'h08: RD = 32'b00000000101000000000000100000011;
			8'h0C: RD = 32'b00000000001000000000010110100011;
			8'h10: RD = 32'b00000000101100000000000110000011;
			8'h14: RD = 32'b00000000001100000000011000100011;
			8'h18: RD = 32'b00000000110000000000001000000011;
			default: RD = 32'b000000_00000_00000_00000_00000_000000;
		endcase
	end
endmodule 
